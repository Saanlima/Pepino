`timescale 1ns / 1ps
// N.Wirth  10.10.2012
module MouseX(
  input clk, enable,
  input [6:0] in,
  output [27:0] out);

  reg x00, x01, x10, x11, y00, y01, y10, y11;
  reg ML, MM, MR;  // keys
  reg [9:0] x, y;  // counters

  wire xup, xdn, yup, ydn;

  assign xup = ~x00&~x01&~x10&x11 | ~x00&x01&x10&x11 | x00&~x01&~x10&~x11 | x00&x01&x10&~x11;
  assign yup = ~y00&~y01&~y10&y11 | ~y00&y01&y10&y11 | y00&~y01&~y10&~y11 | y00&y01&y10&~y11;
  assign xdn = ~x00&~x01&x10&~x11 | ~x00&x01&~x10&~x11 | x00&~x01&x10&x11 | x00&x01&~x10&x11;
  assign ydn = ~y00&~y01&y10&~y11 | ~y00&y01&~y10&~y11 | y00&~y01&y10&y11 | y00&y01&~y10&y11;
  assign out = {1'b0, ML, MM, MR, 2'b0, y, 2'b0, x};
  
  always @ (posedge clk)
    if (enable) begin
      x00 <= in[3]; x01 <= x00; x10 <= in[2]; x11 <= x10;
      y00 <= in[1]; y01 <= y00; y10 <= in[0]; y11 <= y10;
      MR <= ~in[4]; MM <= ~in[5]; ML <= ~in[6];
      x <= xup ? x+1 : xdn ? x-1 : x; 
      y <= yup ? y+1 : ydn ? y-1 : y;
    end
endmodule

